library verilog;
use verilog.vl_types.all;
entity tb_trafficLight is
end tb_trafficLight;
